`timescale 1ns / 1ps

module memory(

    );
endmodule
